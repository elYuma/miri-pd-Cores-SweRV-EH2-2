// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by bscuser on Sat Jan 15 08:53:45 CET 2022
//
// cmd:    swerv -target=default -set=build_axi4 
//

`include "common_defines.vh"
`undef RV_ASSERT_ON
`undef TEC_RV_ICG
`define RV_PHYSICAL 1
